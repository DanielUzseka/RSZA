`ifndef macros_vh
`define macros_vh

`define addrWidth 32
`define dataWidth 32

`endif
