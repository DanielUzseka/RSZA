`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:28:52 04/27/2017 
// Design Name: 
// Module Name:    mod_apb 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module mod_apb(
    input clk,
    input reset,
    input [0:0] addr,
    input [0:0] pwdata,
    input pwrite,
    input psel,
    input penable,
    output [0:0] prdata
    );


endmodule
